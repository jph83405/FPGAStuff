module notGate ( A, B);
  input wire A;
  output wire B;
  assign B=!A;
endmodule // Not gate
